initial begin
    mem[0] = 32'h000002b7;
    mem[1] = 32'h04028293;
    mem[2] = 32'h12345337;
    mem[3] = 32'h6783031b;
    mem[4] = 32'h0062a023;
    mem[5] = 32'h000002b7;
    mem[6] = 32'h04428293;
    mem[7] = 32'h12345337;
    mem[8] = 32'h6783031b;
    mem[9] = 32'h0062a023;
    mem[10] = 32'h000002b7;
    mem[11] = 32'h04828293;
    mem[12] = 32'h12345337;
    mem[13] = 32'h6783031b;
    mem[14] = 32'h0062a023;
    mem[15] = 32'h000002b7;
    mem[16] = 32'h04c28293;
    mem[17] = 32'h12345337;
    mem[18] = 32'h6783031b;
    mem[19] = 32'h0062a023;
    mem[20] = 32'h000002b7;
    mem[21] = 32'h05028293;
    mem[22] = 32'h12345337;
    mem[23] = 32'h6783031b;
    mem[24] = 32'h0062a023;
    mem[25] = 32'h00a00893;
    mem[26] = 32'h00000073;
end