//TO DO
class uart_test extends uvm_test;
    function new();
        
    endfunction //new()
endclass //uart_test extends uvm_test