module top();
    `include "top.vh"
endmodule