//TO DO
class uart_scoreboard extends uvm_scoreboard;
    function new();
        
    endfunction //new()
endclass //uart_scoreboard extends uvm_scoreboard