//TRANSACTION CYCLE:
//1. Start new transaction
//2. Apply control signals
//3. Start transmitter and receiver
//4. Wait for transaction to complete (tx_done and rx_done)
//5. Complete transaction
//6. Repeat