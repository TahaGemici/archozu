// Bootloader code

initial begin
    mem[  0] = 32'h00_00_00_00;
    mem[  1] = 32'h00_00_00_00;
    mem[  2] = 32'h00_00_00_00;
    mem[  3] = 32'h00_00_00_00;
    mem[  4] = 32'h00_00_00_00;
    mem[  5] = 32'h00_00_00_00;
    mem[  6] = 32'h00_00_00_00;
    mem[  7] = 32'h00_00_00_00;
    mem[  8] = 32'h00_00_00_00;
    mem[  9] = 32'h00_00_00_00;
    mem[ 10] = 32'h00_00_00_00;
    mem[ 11] = 32'h00_00_00_00;
    mem[ 12] = 32'h00_00_00_00;
    mem[ 13] = 32'h00_00_00_00;
    mem[ 14] = 32'h00_00_00_00;
    mem[ 15] = 32'h00_00_00_00;
    mem[ 16] = 32'h00_00_00_00;
    mem[ 17] = 32'h00_00_00_00;
    mem[ 18] = 32'h00_00_00_00;
    mem[ 19] = 32'h00_00_00_00;
    mem[ 20] = 32'h00_00_00_00;
    mem[ 21] = 32'h00_00_00_00;
    mem[ 22] = 32'h00_00_00_00;
    mem[ 23] = 32'h00_00_00_00;
    mem[ 24] = 32'h00_00_00_00;
    mem[ 25] = 32'h00_00_00_00;
    mem[ 26] = 32'h00_00_00_00;
    mem[ 27] = 32'h00_00_00_00;
    mem[ 28] = 32'h00_00_00_00;
    mem[ 29] = 32'h00_00_00_00;
    mem[ 30] = 32'h00_00_00_00;
    mem[ 31] = 32'h00_00_00_00;
    mem[ 32] = 32'h00_00_00_00;
    mem[ 33] = 32'h00_00_00_00;
    mem[ 34] = 32'h00_00_00_00;
    mem[ 35] = 32'h00_00_00_00;
    mem[ 36] = 32'h00_00_00_00;
    mem[ 37] = 32'h00_00_00_00;
    mem[ 38] = 32'h00_00_00_00;
    mem[ 39] = 32'h00_00_00_00;
    mem[ 40] = 32'h00_00_00_00;
    mem[ 41] = 32'h00_00_00_00;
    mem[ 42] = 32'h00_00_00_00;
    mem[ 43] = 32'h00_00_00_00;
    mem[ 44] = 32'h00_00_00_00;
    mem[ 45] = 32'h00_00_00_00;
    mem[ 46] = 32'h00_00_00_00;
    mem[ 47] = 32'h00_00_00_00;
    mem[ 48] = 32'h00_00_00_00;
    mem[ 49] = 32'h00_00_00_00;
    mem[ 50] = 32'h00_00_00_00;
    mem[ 51] = 32'h00_00_00_00;
    mem[ 52] = 32'h00_00_00_00;
    mem[ 53] = 32'h00_00_00_00;
    mem[ 54] = 32'h00_00_00_00;
    mem[ 55] = 32'h00_00_00_00;
    mem[ 56] = 32'h00_00_00_00;
    mem[ 57] = 32'h00_00_00_00;
    mem[ 58] = 32'h00_00_00_00;
    mem[ 59] = 32'h00_00_00_00;
    mem[ 60] = 32'h00_00_00_00;
    mem[ 61] = 32'h00_00_00_00;
    mem[ 62] = 32'h00_00_00_00;
    mem[ 63] = 32'h00_00_00_00;
    mem[ 64] = 32'h00_00_00_00;
    mem[ 65] = 32'h00_00_00_00;
    mem[ 66] = 32'h00_00_00_00;
    mem[ 67] = 32'h00_00_00_00;
    mem[ 68] = 32'h00_00_00_00;
    mem[ 69] = 32'h00_00_00_00;
    mem[ 70] = 32'h00_00_00_00;
    mem[ 71] = 32'h00_00_00_00;
    mem[ 72] = 32'h00_00_00_00;
    mem[ 73] = 32'h00_00_00_00;
    mem[ 74] = 32'h00_00_00_00;
    mem[ 75] = 32'h00_00_00_00;
    mem[ 76] = 32'h00_00_00_00;
    mem[ 77] = 32'h00_00_00_00;
    mem[ 78] = 32'h00_00_00_00;
    mem[ 79] = 32'h00_00_00_00;
    mem[ 80] = 32'h00_00_00_00;
    mem[ 81] = 32'h00_00_00_00;
    mem[ 82] = 32'h00_00_00_00;
    mem[ 83] = 32'h00_00_00_00;
    mem[ 84] = 32'h00_00_00_00;
    mem[ 85] = 32'h00_00_00_00;
    mem[ 86] = 32'h00_00_00_00;
    mem[ 87] = 32'h00_00_00_00;
    mem[ 88] = 32'h00_00_00_00;
    mem[ 89] = 32'h00_00_00_00;
    mem[ 90] = 32'h00_00_00_00;
    mem[ 91] = 32'h00_00_00_00;
    mem[ 92] = 32'h00_00_00_00;
    mem[ 93] = 32'h00_00_00_00;
    mem[ 94] = 32'h00_00_00_00;
    mem[ 95] = 32'h00_00_00_00;
    mem[ 96] = 32'h00_00_00_00;
    mem[ 97] = 32'h00_00_00_00;
    mem[ 98] = 32'h00_00_00_00;
    mem[ 99] = 32'h00_00_00_00;
    mem[100] = 32'h00_00_00_00;
    mem[101] = 32'h00_00_00_00;
    mem[102] = 32'h00_00_00_00;
    mem[103] = 32'h00_00_00_00;
    mem[104] = 32'h00_00_00_00;
    mem[105] = 32'h00_00_00_00;
    mem[106] = 32'h00_00_00_00;
    mem[107] = 32'h00_00_00_00;
    mem[108] = 32'h00_00_00_00;
    mem[109] = 32'h00_00_00_00;
    mem[110] = 32'h00_00_00_00;
    mem[111] = 32'h00_00_00_00;
    mem[112] = 32'h00_00_00_00;
    mem[113] = 32'h00_00_00_00;
    mem[114] = 32'h00_00_00_00;
    mem[115] = 32'h00_00_00_00;
    mem[116] = 32'h00_00_00_00;
    mem[117] = 32'h00_00_00_00;
    mem[118] = 32'h00_00_00_00;
    mem[119] = 32'h00_00_00_00;
    mem[120] = 32'h00_00_00_00;
    mem[121] = 32'h00_00_00_00;
    mem[122] = 32'h00_00_00_00;
    mem[123] = 32'h00_00_00_00;
    mem[124] = 32'h00_00_00_00;
    mem[125] = 32'h00_00_00_00;
    mem[126] = 32'h00_00_00_00;
    mem[127] = 32'h00_00_00_00;
end