interface uart_interface;
    //TO DO
endinterface //uart_interface//TO DO